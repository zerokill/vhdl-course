-- Test Bench voor opdracht 3
-- Datum : 18 Mei 2007
-- E.G. van den Bor
-- Hogeschool Utrecht
--
-- In deze testbench worden een aantal constanten aan ingang A en B
-- gegeven.
-- Bij alle combinaties van de Code (deel van een ALU instructie)
-- wordt het resultaat van de aangeboden constanten gecontroleerd.
-- Deze testbench bestaat uit vijf processen
-- Dit zijn :
-- Stim_A en Stim_B : hierin worden de constanten gekoppeld aan ingang A en B
-- Stim_code : Hierin wordt de Code voor iedere bewerking bepaald
-- Expected : Hierin wordt de verwachtw waarde berekend
-- Controle : controleert of de uitgang overeen komt met de verwachte waarde
-- de vijf processen lopen parallel (concurrent).
-- Na iedere 10 ns is er een nieuw resultaat bekend.
-- De controle vindt plaats net voordat een nieuwe waarde wordt aangboden
-- Namelijk na 9 ns Zodat het uitgangssignaal stabiel is.

entity ALU_TB is
end;

library IEEE;
use IEEE.Std_logic_1164.all;
use IEEE.Numeric_Std.all;

architecture Bench of ALU_TB is

  constant OP_SIZE       : POSITIVE := 4; -- breedte van de opcode

  -- Signalen die aan de ALU file worden verbonden
  -- ingangen van de ALU  
  signal A, B: std_logic_vector(7 downto 0) := (others => '0');
  signal Code: std_logic_vector(OP_SIZE-1 downto 0);
  -- uitgangen van de ALU
  signal Cout, Equal : Std_logic;
  signal F: std_logic_vector(7 downto 0);

  
  -- De onderstaande constanten worden als testwaarden
  -- gebruikt van zowel ingang A als B bij iedere mogelijke
  -- bewerking
  constant Value0: Std_logic_vector := "00000000";
  constant Value1: Std_logic_vector := "00000001";
  constant Value2: Std_logic_vector := "00000011";
  constant Value3: Std_logic_vector := "00001000";
  constant Value4: Std_logic_vector := "00001111";
  constant Value5: Std_logic_vector := "10000000";
  constant Value6: Std_logic_vector := "11111000";
  constant Value7: Std_logic_vector := "11111111";

  constant NUM_TESTCONST    : POSITIVE := 8; -- aantal testconstanten
  constant NUM_OPCODES      : POSITIVE := 2 ** OP_SIZE; -- aantal opcodes
  constant NUM_TOT_VECTORS  : POSITIVE := NUM_TESTCONST * NUM_TESTCONST * NUM_OPCODES;
  -- totaal aantal testvectoren
  
  -- Vertragingstijden 
  constant OP_DELAY : TIME := 10 ns;
  constant  A_DELAY : TIME := NUM_OPCODES * OP_DELAY;
  constant  B_DELAY : TIME := NUM_TESTCONST * A_DELAY;

  -- Verwachte resultaten en fouttellers
  signal Verwacht : Std_logic_vector(1 to 10);   -- hierin komen de 
  -- verwachte resultaten
  constant DONT_CARE : Std_logic_vector(7 downto 0) := "--------";

  signal     F_fout_teller : NATURAL := 0;
  signal  Cout_fout_teller : NATURAL := 0;
  signal Equal_fout_teller : NATURAL := 0;

  signal     F_OK : BOOLEAN := TRUE;
  signal  Cout_OK : BOOLEAN := TRUE;
  signal Equal_OK : BOOLEAN := TRUE;

begin
-- Koppel eerste de testbench file aan de ALU file
  UUT: entity work.ALU port map ( 
					A     => A,
               B     => B,
               Code  => Code,
               F     => F,
               Cout  => Cout,
               Equal => Equal);

  -- Koppel aan ingang B steeds een testconstante
  Stim_B: process
  begin
    B <= Value0;
    wait for B_DELAY;
    B <= Value1;
    wait for B_DELAY;
    B <= Value2;
    wait for B_DELAY;
    B <= Value3;
    wait for B_DELAY;
    B <= Value4;
    wait for B_DELAY;
    B <= Value5;
    wait for B_DELAY;
    B <= Value6;
    wait for B_DELAY;
    B <= Value7;
    wait for B_DELAY;
    wait;
  end process Stim_B;

  -- Koppel aan ingang A steeds een testconstante
  -- terwijl ingang B tijdelijk gelijk blijft
  Stim_A: process
  begin
    for I in 1 to NUM_TESTCONST loop
      A <= Value0;
      wait for A_DELAY;
      A <= Value1;
      wait for A_DELAY;
      A <= Value2;
      wait for A_DELAY;
      A <= Value3;
      wait for A_DELAY;
      A <= Value4;
      wait for A_DELAY;
      A <= Value5;
      wait for A_DELAY;
      A <= Value6;
      wait for A_DELAY;
      A <= Value7;
      wait for A_DELAY;
    end loop;
    wait;
  end process Stim_A;

  -- Geef de Opcode bij alle mogelijke combinaties van A en B
  -- inclusief de niet gebruikte opcodes
  
  Stim_Code: process
  begin
    for I in 1 to NUM_TESTCONST * NUM_TESTCONST loop
      for J in 0 to NUM_OPCODES-1 loop
        Code <= Std_logic_vector(To_unsigned(J,4));
        wait for OP_DELAY;
      end loop;
    end loop;
    wait;
  end process Stim_Code;

  -- Geef de verwachte waarden en plaats die in het signal "Verwacht".
  Expected: process
  begin
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "1000000100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "1000011100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000010"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "0000000110"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111000010"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111010"; wait for OP_DELAY;
    Verwacht <= "0111111100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000001001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000000101"; wait for OP_DELAY;
    Verwacht <= "0000000101"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "0000001001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000001001"; wait for OP_DELAY;
    Verwacht <= "1000000001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "1111111010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "1000000100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000100100"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "1111100110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000111000"; wait for OP_DELAY;
    Verwacht <= "1111001010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "1000011100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000000110"; wait for OP_DELAY;
    Verwacht <= "0111111110"; wait for OP_DELAY;
    Verwacht <= "1000000100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000010"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "0000000110"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111100110"; wait for OP_DELAY;
    Verwacht <= "1111011110"; wait for OP_DELAY;
    Verwacht <= "0000100100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111000010"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111010"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111010"; wait for OP_DELAY;
    Verwacht <= "0111111100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "1111111010"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000011001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000001101"; wait for OP_DELAY;
    Verwacht <= "0000001101"; wait for OP_DELAY;
    Verwacht <= "1111110111"; wait for OP_DELAY;
    Verwacht <= "1111110111"; wait for OP_DELAY;
    Verwacht <= "0000011001"; wait for OP_DELAY;
    Verwacht <= "0000000101"; wait for OP_DELAY;
    Verwacht <= "0000011001"; wait for OP_DELAY;
    Verwacht <= "1000000101"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "0000101100"; wait for OP_DELAY;
    Verwacht <= "0000010100"; wait for OP_DELAY;
    Verwacht <= "1111101110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0001001000"; wait for OP_DELAY;
    Verwacht <= "0000110000"; wait for OP_DELAY;
    Verwacht <= "1111010010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "1000011100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000001110"; wait for OP_DELAY;
    Verwacht <= "0111110110"; wait for OP_DELAY;
    Verwacht <= "1000001100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "0000000010"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "0000000110"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111101110"; wait for OP_DELAY;
    Verwacht <= "1111010110"; wait for OP_DELAY;
    Verwacht <= "0000101100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "1111000010"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "1111110010"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "1111111010"; wait for OP_DELAY;
    Verwacht <= "0111111100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000100100"; wait for OP_DELAY;
    Verwacht <= "1111100110"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000101100"; wait for OP_DELAY;
    Verwacht <= "1111101110"; wait for OP_DELAY;
    Verwacht <= "0000010100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "1000000100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0001000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000100001"; wait for OP_DELAY;
    Verwacht <= "0000100001"; wait for OP_DELAY;
    Verwacht <= "1111100011"; wait for OP_DELAY;
    Verwacht <= "1111100011"; wait for OP_DELAY;
    Verwacht <= "0001000001"; wait for OP_DELAY;
    Verwacht <= "0000010001"; wait for OP_DELAY;
    Verwacht <= "0001000001"; wait for OP_DELAY;
    Verwacht <= "0000010001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "0001011100"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "1111100110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "1000011100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000100010"; wait for OP_DELAY;
    Verwacht <= "0111100010"; wait for OP_DELAY;
    Verwacht <= "1000100000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000000010"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "0000000110"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111000010"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1111000010"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "1111011110"; wait for OP_DELAY;
    Verwacht <= "0000100100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1111111010"; wait for OP_DELAY;
    Verwacht <= "0111111100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "1111001010"; wait for OP_DELAY;
    Verwacht <= "0000111000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0001001000"; wait for OP_DELAY;
    Verwacht <= "1111010010"; wait for OP_DELAY;
    Verwacht <= "0000110000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "1000000100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0001011100"; wait for OP_DELAY;
    Verwacht <= "1111100110"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0001111001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000111101"; wait for OP_DELAY;
    Verwacht <= "0000111101"; wait for OP_DELAY;
    Verwacht <= "1111000111"; wait for OP_DELAY;
    Verwacht <= "1111000111"; wait for OP_DELAY;
    Verwacht <= "0001111001"; wait for OP_DELAY;
    Verwacht <= "0000011101"; wait for OP_DELAY;
    Verwacht <= "0001111001"; wait for OP_DELAY;
    Verwacht <= "1000011101"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "1000111110"; wait for OP_DELAY;
    Verwacht <= "0111000110"; wait for OP_DELAY;
    Verwacht <= "1000111100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0000000010"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "0000000110"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "1110100110"; wait for OP_DELAY;
    Verwacht <= "0001011100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "1111000010"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000111000"; wait for OP_DELAY;
    Verwacht <= "1111000010"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "1111111010"; wait for OP_DELAY;
    Verwacht <= "0111111100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000000110"; wait for OP_DELAY;
    Verwacht <= "1000000100"; wait for OP_DELAY;
    Verwacht <= "0111111110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000001110"; wait for OP_DELAY;
    Verwacht <= "1000001100"; wait for OP_DELAY;
    Verwacht <= "0111110110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "1000000100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000100010"; wait for OP_DELAY;
    Verwacht <= "1000100000"; wait for OP_DELAY;
    Verwacht <= "0111100010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000111110"; wait for OP_DELAY;
    Verwacht <= "1000111100"; wait for OP_DELAY;
    Verwacht <= "0111000110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "1000011100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000011"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "1000000011"; wait for OP_DELAY;
    Verwacht <= "1000000011"; wait for OP_DELAY;
    Verwacht <= "1000000001"; wait for OP_DELAY;
    Verwacht <= "1000000001"; wait for OP_DELAY;
    Verwacht <= "0000000011"; wait for OP_DELAY;
    Verwacht <= "0100000001"; wait for OP_DELAY;
    Verwacht <= "0000000111"; wait for OP_DELAY;
    Verwacht <= "0100000001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "0111100010"; wait for OP_DELAY;
    Verwacht <= "0111100000"; wait for OP_DELAY;
    Verwacht <= "1000100010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "1111000010"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0111111110"; wait for OP_DELAY;
    Verwacht <= "0111111100"; wait for OP_DELAY;
    Verwacht <= "1000000110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "1111111010"; wait for OP_DELAY;
    Verwacht <= "0111111100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111100110"; wait for OP_DELAY;
    Verwacht <= "0000100100"; wait for OP_DELAY;
    Verwacht <= "1111011110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111101110"; wait for OP_DELAY;
    Verwacht <= "0000101100"; wait for OP_DELAY;
    Verwacht <= "1111010110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "1000000100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "1111000010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "0001011100"; wait for OP_DELAY;
    Verwacht <= "1110100110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "1000011100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0111100010"; wait for OP_DELAY;
    Verwacht <= "1000100010"; wait for OP_DELAY;
    Verwacht <= "0111100000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000000010"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "0000000110"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111000011"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "1111100011"; wait for OP_DELAY;
    Verwacht <= "1111100011"; wait for OP_DELAY;
    Verwacht <= "0000100001"; wait for OP_DELAY;
    Verwacht <= "0000100001"; wait for OP_DELAY;
    Verwacht <= "1111000011"; wait for OP_DELAY;
    Verwacht <= "0111110001"; wait for OP_DELAY;
    Verwacht <= "1111000111"; wait for OP_DELAY;
    Verwacht <= "0111110001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "1111011110"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "1111100110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111111010"; wait for OP_DELAY;
    Verwacht <= "0111111100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "1111111010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000001000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "1111110010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000001100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111110110"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000011000"; wait for OP_DELAY;
    Verwacht <= "1000000100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "0000100100"; wait for OP_DELAY;
    Verwacht <= "1111011110"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "0000010000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000111000"; wait for OP_DELAY;
    Verwacht <= "0001000000"; wait for OP_DELAY;
    Verwacht <= "1111000010"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000111100"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "0001111000"; wait for OP_DELAY;
    Verwacht <= "1000011100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0111111110"; wait for OP_DELAY;
    Verwacht <= "1000000110"; wait for OP_DELAY;
    Verwacht <= "0111111100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1000000010"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1000000000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "0000000010"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "0000000110"; wait for OP_DELAY;
    Verwacht <= "0100000000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111011110"; wait for OP_DELAY;
    Verwacht <= "1111100110"; wait for OP_DELAY;
    Verwacht <= "0000011100"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "1111100010"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "0000100000"; wait for OP_DELAY;
    Verwacht <= "0000000100"; wait for OP_DELAY;
    Verwacht <= "1111000010"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "1111000110"; wait for OP_DELAY;
    Verwacht <= "0111110000"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "---------0"; wait for OP_DELAY;
    Verwacht <= "0000000000"; wait for OP_DELAY;
    Verwacht <= "1111111110"; wait for OP_DELAY;
    Verwacht <= "1111111011"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "0000000101"; wait for OP_DELAY;
    Verwacht <= "0000000101"; wait for OP_DELAY;
    Verwacht <= "1111111011"; wait for OP_DELAY;
    Verwacht <= "0111111101"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    Verwacht <= "1111111101"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "---------1"; wait for OP_DELAY;
    Verwacht <= "0000000001"; wait for OP_DELAY;
    Verwacht <= "1111111111"; wait for OP_DELAY;
    wait;
  end process Expected;

  -- Dit process controleert of de verwachte resultaten 
  -- overeenstemmen met die uit de VHDL file.
  -- Bij verwachte don't care waarde ('_') wordt de uitgang van de 
  -- VHDL file gegegeerd.
  Controle : process
  begin
    wait for OP_DELAY - 1 NS;
    for I in 1 to NUM_TOT_VECTORS loop
      -- Hieronder staat de controle van uitgang F
      if ( Verwacht(1 to 8) /= DONT_CARE ) and ( F /= Verwacht(1 to 8) ) then
        F_OK              <= FALSE;
        F_fout_teller     <= F_fout_teller + 1;
      end if;
      -- Hieronder staat de controle Carry out
      if ( Verwacht(9) /= '-' ) and ( Cout /= Verwacht(9) ) then
        Cout_OK           <= FALSE;
        Cout_fout_teller  <= Cout_fout_teller + 1;
      end if;
      -- Hieronder staat de controle equal uitgang
      if ( Verwacht(10) /= '-' ) and ( Equal /= Verwacht(10) ) then
        Equal_OK          <= FALSE;
        Equal_fout_teller <= Equal_fout_teller + 1;
      end if;
      wait for OP_DELAY;
    end loop;
    wait;
  end process Controle;

end architecture Bench;
